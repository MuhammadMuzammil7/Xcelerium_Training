// Layered Testbench of Shift Register:
// Shift Register Transaction Class
class shift_reg_transaction #(parameter N = 8);
    rand bit shift_en;
    rand bit dir;
    rand bit d_in;
    bit [N-1:0] q_out;
    
    constraint valid_c {
        shift_en dist {1 := 80, 0 := 20};
        dir dist {0 := 50, 1 := 50};
    }
    
    function void display(string tag = "");
        $display("[%0t] %s: shift_en=%0b, dir=%0s, d_in=%0b, q_out=%0h", 
                 $time, tag, shift_en, dir ? "RIGHT" : "LEFT", d_in, q_out);
    endfunction
endclass

// Shift Register Generator Class
class shift_reg_generator #(parameter N = 8);
    mailbox #(shift_reg_transaction#(N)) gen2drv;
    int num_trans;
    
    function new(mailbox #(shift_reg_transaction#(N)) g2d, int n = 100);
        this.gen2drv = g2d;
        this.num_trans = n;
    endfunction
    
    task run();
        shift_reg_transaction#(N) trans;
        repeat(num_trans) begin
            trans = new();
            assert(trans.randomize()) else $fatal("Randomization failed");
            gen2drv.put(trans);
        end
    endtask
endclass

// Shift Register Driver Class
class shift_reg_driver #(parameter N = 8);
    virtual shift_reg_if#(N) vif;
    mailbox #(shift_reg_transaction#(N)) gen2drv;
    
    function new(virtual shift_reg_if#(N) vif, mailbox #(shift_reg_transaction#(N)) g2d);
        this.vif = vif;
        this.gen2drv = g2d;
    endfunction
    
    task reset();
        vif.rst_n <= 0;
        vif.shift_en <= 0;
        vif.dir <= 0;
        vif.d_in <= 0;
        repeat(2) @(posedge vif.clk);
        vif.rst_n <= 1;
        @(posedge vif.clk);
    endtask
    
    task run();
        shift_reg_transaction#(N) trans;
        forever begin
            gen2drv.get(trans);
            @(posedge vif.clk);
            vif.shift_en <= trans.shift_en;
            vif.dir <= trans.dir;
            vif.d_in <= trans.d_in;
            trans.display("DRIVER");
        end
    endtask
endclass

// Shift Register Monitor Class
class shift_reg_monitor #(parameter N = 8);
    virtual shift_reg_if#(N) vif;
    mailbox #(shift_reg_transaction#(N)) mon2scb;
    
    function new(virtual shift_reg_if#(N) vif, mailbox #(shift_reg_transaction#(N)) m2s);
        this.vif = vif;
        this.mon2scb = m2s;
    endfunction
    
    task run();
        shift_reg_transaction#(N) trans;
        forever begin
            @(posedge vif.clk);
            trans = new();
            trans.shift_en = vif.shift_en;
            trans.dir = vif.dir;
            trans.d_in = vif.d_in;
            trans.q_out = vif.q_out;
            mon2scb.put(trans);
            trans.display("MONITOR");
        end
    endtask
endclass

// Shift Register Scoreboard Class
class shift_reg_scoreboard #(parameter N = 8);
    mailbox #(shift_reg_transaction#(N)) mon2scb;
    bit [N-1:0] expected_q;
    int pass_count, fail_count;
    
    function new(mailbox #(shift_reg_transaction#(N)) m2s);
        this.mon2scb = m2s;
        this.expected_q = 0;
        this.pass_count = 0;
        this.fail_count = 0;
    endfunction
    
    task run();
        shift_reg_transaction#(N) trans;
        forever begin
            mon2scb.get(trans);
            
            if (trans.q_out === expected_q) begin
                $display("[%0t] SCOREBOARD PASS: Expected=%0h, Got=%0h", 
                         $time, expected_q, trans.q_out);
                pass_count++;
            end else begin
                $display("[%0t] SCOREBOARD FAIL: Expected=%0h, Got=%0h", 
                         $time, expected_q, trans.q_out);
                fail_count++;
            end
            
            // Update expected output
            if (trans.shift_en) begin
                if (trans.dir) // Right shift
                    expected_q = {trans.d_in, expected_q[N-1:1]};
                else // Left shift
                    expected_q = {expected_q[N-2:0], trans.d_in};
            end
        end
    endtask
    
    function void report();
        $display("\n========== SCOREBOARD REPORT ==========");
        $display("Total Passed: %0d", pass_count);
        $display("Total Failed: %0d", fail_count);
        $display("=======================================\n");
    endfunction
endclass

// Shift Register Environment Class
class shift_reg_environment #(parameter N = 8);
    shift_reg_generator#(N) gen;
    shift_reg_driver#(N) drv;
    shift_reg_monitor#(N) mon;
    shift_reg_scoreboard#(N) scb;
    
    mailbox #(shift_reg_transaction#(N)) gen2drv;
    mailbox #(shift_reg_transaction#(N)) mon2scb;
    
    virtual shift_reg_if#(N) vif;
    
    function new(virtual shift_reg_if#(N) vif);
        this.vif = vif;
        gen2drv = new();
        mon2scb = new();
        
        gen = new(gen2drv, 100);
        drv = new(vif, gen2drv);
        mon = new(vif, mon2scb);
        scb = new(mon2scb);
    endfunction
    
    task run();
        fork
            drv.reset();
            #100 gen.run();
            drv.run();
            mon.run();
            scb.run();
        join_any
    endtask
    
    function void report();
        scb.report();
    endfunction
endclass

// Shift Register Interface
interface shift_reg_if #(parameter N = 8)(input logic clk);
    logic rst_n;
    logic shift_en;
    logic dir;
    logic d_in;
    logic [N-1:0] q_out;
endinterface

// Shift Register Testbench Top
module shift_reg_tb;
    parameter N = 8;
    logic clk;
    
    shift_reg_if#(N) sif(clk);
    
    shift_reg#(N) dut (
        .clk(sif.clk),
        .rst_n(sif.rst_n),
        .shift_en(sif.shift_en),
        .dir(sif.dir),
        .d_in(sif.d_in),
        .q_out(sif.q_out)
    );
    
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end
    
    shift_reg_environment#(N) env;
    
    initial begin
        env = new(sif);
        env.run();
        #2000;
        env.report();
        $finish;
    end

    // Dump waveforms
    initial begin
        $dumpfile("shift_reg.vcd");
        $dumpvars(0, shift_reg_tb_layered);
    end
endmodule